/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-22 20:52:35 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-23 12:23:20
 */

 // parameter define
 `define true   1'b1
 `define false  1'b0


 