/home/dracacys/ics2023/npc/naive_cpu/vsrc/INST_MEM.sv