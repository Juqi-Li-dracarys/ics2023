/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-21 15:56:01 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-21 16:54:07
 */

// parameter define
 `define true   1'b1
 `define false  1'b0

// parameter define
`define PC_RST 32'h80000000
`define NOP    32'h00000013

// master state
`define  idle       1'b0
`define  wait_ready 1'b1


