/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-19 13:23:33 
 * @Last Modified by:   Juqi Li @ NJU 
 * @Last Modified time: 2024-02-19 13:23:33 
 */

 `include "IDU_DEFINES_ysyx23060136.sv"


 