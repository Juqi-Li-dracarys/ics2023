/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-27 16:42:25 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-27 16:42:45
 */



module WB_TOP_ysyx23060136 (
    
);
    
endmodule


