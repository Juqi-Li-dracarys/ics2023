/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-17 15:02:46 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-21 16:56:15
 */


// parameter define
 `define true   'b1
 `define false  'b0

// csr idx 
`define  mstatus  2'h0 
`define  mtvec    2'h1
`define  mepc     2'h2
`define  mcause   2'h3

        
