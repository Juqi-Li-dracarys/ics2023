/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-24 17:15:34 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-24 17:16:15
 */

 module MEM_FORWARD_ysyx23060136 (

 );
    
endmodule



 
