/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-28 13:07:41 
 * @Last Modified by:   Juqi Li @ NJU 
 * @Last Modified time: 2024-02-28 13:07:41 
 */


 module MEM_TOP_ysyx23060136 (

 );
    
endmodule

