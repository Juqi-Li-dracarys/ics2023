/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-24 21:16:59 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-24 21:20:00
 */

 module MEM_SRAM_ysyx23060136 (

 );
    
endmodule



