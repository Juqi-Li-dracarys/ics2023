/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-24 17:17:00 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-24 17:17:20
 */

 module MEM_TOP_ysyx23060136 (

 );
    
endmodule

