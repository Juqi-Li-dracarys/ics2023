/home/dracacys/ics2023/npc/naive_cpu/vsrc/CPU_TOP.sv