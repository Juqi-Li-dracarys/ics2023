
`include "../include/interface_ysyx23060136.svh"


module SRAM_ysyx23060136(

);

endmodule

