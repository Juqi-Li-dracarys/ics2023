/home/dracacys/ics2023/npc/naive_cpu/vsrc/ALU.sv