/home/dracacys/ics2023/npc/naive_cpu/vsrc/CRTL_GEN.sv