/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-15 23:40:06 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-17 15:04:14
 */

`include "IDU_DEFINES_ysyx23060136.sv"

///////////////////////////////////////////////

module IDU_IMM_GEN_ysyx_23060136(
        input         [31 : 7]   inst,
        input         [2 : 0]    opcode,   // 指令类型
        output logic  [31 : 0]   imm
    );

    always_comb begin
        unique case(opcode)
            `I_type:                                                                          // I type
                imm = {{20{inst[31]}}, inst[31 : 20]};
            `S_type:                                                                          // S type
                imm = {{20{inst[31]}}, inst[31 : 25], inst[11 : 7]};
            `B_type:                                                                          // B type
                imm = {{20{inst[31]}}, inst[7], inst[30 : 25], inst[11 : 8], 1'b0};
            `U_type:                                                                          // U type
                imm = {inst[31 : 12], 12'b0};
            `J_type:                                                                          // J type
                imm = {{12{inst[31]}}, inst[19 : 12], inst[20], inst[30 : 21], 1'b0};
            default:
                imm = 32'b0;                                                                  // R-type
        endcase
    end

endmodule



