/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-04-18 16:28:13 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-04-18 16:29:47
 */


module  ysyx_23060136_MEM_AXI(
   
);
    
endmodule



