/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-16 13:50:37 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-16 13:53:16
 */


// parameter define
 `define true   1'b1
 `define false  1'b0

// parameter define
`define PC_RST 32'h80000000

// master state
`define  idle       1'b0
`define  wait_ready 1'b1

        
