/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-24 01:40:32 
 * @Last Modified by:   Juqi Li @ NJU 
 * @Last Modified time: 2024-02-24 01:40:32 
 */
module moduleName (
    ports
);
    
endmodule