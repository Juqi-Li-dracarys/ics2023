/home/dracacys/ics2023/npc/naive_cpu/vsrc/PC_SEL.sv