/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-24 17:17:47 
 * @Last Modified by:   Juqi Li @ NJU 
 * @Last Modified time: 2024-02-24 17:17:47 
 */

