/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-01-14 09:07:03 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-01-14 10:36:45
 */


module CPU_TOP #(parameter PC_RST = 32'h80000000) (
    input                      clk, rst,
    output      [31: 0]        pc_cur, inst,
    output                     reg_signal,
    output                     inst_signal
);

// TO DO

endmodule


