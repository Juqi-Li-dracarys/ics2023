/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-17 15:02:46 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-17 15:05:25
 */


// parameter define
 `define true   1'b1
 `define false  1'b0

 
// 指令立即数提取

`define   I_type   3'b000
`define   S_type   3'b010
`define   B_type   3'b011
`define   U_type   3'b001
`define   J_type   3'b100
`define   R_type   3'b111

// something wrong
`define   N_type   3'b101
        
