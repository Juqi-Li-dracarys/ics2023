/*
 * @Author: Juqi Li @ NJU 
 * @Date: 2024-02-16 13:50:37 
 * @Last Modified by: Juqi Li @ NJU
 * @Last Modified time: 2024-02-24 23:18:43
 */


// parameter define
 `define true   'b1
 `define false  'b0

// parameter define
`define PC_RST 32'h80000000

// master state
`define  idle       2'h0
`define  busy       2'h1
`define  done       2'h2

        
